/*
CS 274
Ursinus College

@author Michael Cummins
@purpose Implementation control unit
*/

`include "control_unit.v"
`default_nettype none
`timescale 1ns / 1ps

module program();


endmodule